//-------------------------------------------------------------------------------------------------
module ram
//-------------------------------------------------------------------------------------------------
#
(
	parameter KB = 0
)
(
	input  wire                      clock,
	input  wire[$clog2(KB*1024)-1:0] a,
	input  wire[                7:0] d,
	output reg [                7:0] q,
	input  wire                      w
);
//-------------------------------------------------------------------------------------------------

reg[7:0] mem[0:(KB*1024)-1];

always @(posedge clock) if(w) begin mem[a] <= d; q <= d; end else q <= mem[a];

//-------------------------------------------------------------------------------------------------
endmodule
//-------------------------------------------------------------------------------------------------
//-------------------------------------------------------------------------------------------------
module ramm
//-------------------------------------------------------------------------------------------------
#
(
	parameter KB = 0,
	parameter FN = ""
)
(
	input  wire                      clock,
	input  wire[$clog2(KB*1024)-1:0] a,
	input  wire[                7:0] d,
	output reg [                7:0] q,
	input  wire                      w
);
//-------------------------------------------------------------------------------------------------

(* ram_init_file = FN *) reg[7:0] mem[0:(KB*1024)-1];

always @(posedge clock) if(w) begin mem[a] <= d; q <= d; end else q <= mem[a];

//-------------------------------------------------------------------------------------------------
endmodule
//-------------------------------------------------------------------------------------------------
