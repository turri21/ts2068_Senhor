//-------------------------------------------------------------------------------------------------
module romm
//-------------------------------------------------------------------------------------------------
#
(
	parameter KB = 0,
	parameter FN = ""
)
(
	input  wire                      clock,
	input  wire[$clog2(KB*1024)-1:0] a,
	output reg [                7:0] q
);
//-------------------------------------------------------------------------------------------------

(* ram_init_file = FN *) reg[7:0] mem[0:(KB*1024)-1];

reg[7:0] d = 8'hFF;
reg      w = 1'b0;

always @(posedge clock) if(w) begin mem[a] <= d; q <= d; end else q <= mem[a];

//-------------------------------------------------------------------------------------------------
endmodule
//-------------------------------------------------------------------------------------------------
